// $Id: $
// File name:   fifo_RAM.sv
// Created:     4/21/2016
// Author:      Jordan Huffaker
// Lab Section: 337-08
// Version:     1.0  Initial Design Entry
// Description: An abstracted version of RAM as a FIFO.

module fifo_RAM
(
	input wire clk,
	input wire reset,
	input wire write,
	input wire read,
	input wire [31:0] r_data,
	input wire [31:0] w_data,
	output wire empty,
	output wire full
);

	reg []

endmodule
